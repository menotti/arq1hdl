library ieee;
use ieee.std_logic_1164.all;

entity ram is
   generic (
       DATA_WIDTH : natural := 8;
       ADDR_WIDTH : natural := 8);
   port (
       clk: in std_logic;
       addr_a: in natural range 0 to 2**ADDR_WIDTH - 1; 
       addr_b: in natural range 0 to 2**ADDR_WIDTH - 1; 
       data_a: in std_logic_vector((DATA_WIDTH-1) downto 0); 
       data_b: in std_logic_vector((DATA_WIDTH-1) downto 0); 
       we_a: in std_logic := '1';
       we_b: in std_logic := '1';
       q_a: out std_logic_vector((DATA_WIDTH -1) downto 0); 
       q_b: out std_logic_vector((DATA_WIDTH -1) downto 0));
end ram;

architecture rtl of ram is
   -- Build a 2-D array type for the RAM
   subtype word_t is std_logic_vector((DATA_WIDTH-1) downto 0);
   type memory_t is array((2**ADDR_WIDTH - 1) downto 0) of word_t;
   -- Declare the RAM signal.
   shared variable ram : memory_t := (
     0 => "10000000000000000000000000000000",
     1 => "00000000000000000000000000000000",
     2 => "00000000000000000000000000000000",
     3 => "00000000000000000000000000000000",
     4 => "00000000000000000000000000000000",
     5 => "00000000000000000000000000000000",
     6 => "00000000000000000000000000000000",
     7 => "00000000000000000000000000000000",
     8 => "00000000000000000000000000000000",
     9 => "00000000000000000000000000000001",
	  10 => "00011111000110000000000000000000",
    11 => "00000000000000000000000000000000",
    12 => "00000000000000000000000000000000",
    13 => "00000000000000000000000000000000",
    14 => "00000000000000000000000000000000",
    15 => "00000000000000000000000000000000",
    16 => "00000000000000000000000000000000",
    17 => "00000000000000000000000000000000",
    18 => "00000000000000000000000000000000",
    19 => "00000000000000000000000000000001",
	  20 => "00110001100000000000000000000000",
    21 => "00000000000000000000000000000000",
    22 => "00000000000000000000000000000000",
    23 => "00000000000000000000000000000000",
    24 => "00000000000000000000000000000000",
    25 => "00000000000000000000000000000000",
    26 => "00000000000000000000000000000000",
    27 => "00000000000000000000000000000000",
    28 => "00000000000000000000000000000000",
    29 => "00000000000000000000000000000001",
	  30 => "00110001100110000000000000000000",
    31 => "00000000000000000000000000000000",
    32 => "00000000000000000000000000000000",
    33 => "00000000000000000000000000000000",
    34 => "00000000000000000000000000000000",
    35 => "00000000000000000000000000000000",
    36 => "00000000000000000000000000000000",
    37 => "00000000000000000000000000000000",
    38 => "00000000000000000000000000000000",
    39 => "00000000000000000000000000000001",
	  40 => "00110001100110000000000000000000",
    41 => "00000000000000000000000000000000",
    42 => "00000000000000000000000000000000",
    43 => "00000000000000000000000000000000",
    44 => "00000000000000000000000000000000",
    45 => "00000000000000000000000000000000",
    46 => "00000000000000000000000000000000",
    47 => "00000000000000000000000000000000",
    48 => "00000000000000000000000000000000",
    49 => "00000000000000000000000000000001",
	  50 => "00011111000110000000000000000000",
    51 => "00000000000000000000000000000000",
    52 => "00000000000000000000000000000000",
    53 => "00000000000000000000000000000000",
    54 => "00000000000000000000000000000000",
    55 => "00000000000000000000000000000000",
    56 => "00000000000000000000000000000000",
    57 => "00000000000000000000000000000000",
    58 => "00000000000000000000000000000000",
    59 => "00000000000000000000000000000001",
	  60 => "00000000000000000000000000000000",
    61 => "00000000000000000000000000000000",
    62 => "00000000000000000000000000000000",
    63 => "00000000000000000000000000000000",
    64 => "00000000000000000000000000000000",
    65 => "00000000000000000000000000000000",
    66 => "00000000000000000000000000000000",
    67 => "00000000000000000000000000000000",
    68 => "00000000000000000000000000000000",
    69 => "00000000000000000000000000000001",
		others => "10101010101010101010101010101010");
     
   begin

   process(clk)
   begin
   if(rising_edge(clk)) then -- Port B
       if(we_b = '1') then
          ram(addr_b) := data_b;
          -- Read-during-write on the same port returns NEW data
          q_b <= data_b;
       else
          -- Read-during-write on the mixed port returns OLD data
          q_b <= ram(addr_b);
       end if;
   end if;
   end process;

   process(clk)
   begin
   if(rising_edge(clk)) then -- Port A
       if(we_a = '1') then
          ram(addr_a) := data_a;
          -- Read-during-write on the same port returns NEW data
          q_a <= data_a;
       else
          -- Read-during-write on the mixed port returns OLD data
          q_a <= ram(addr_a);
       end if;
   end if;
   end process;
   
end rtl;